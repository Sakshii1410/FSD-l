<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-656.1,86.2,801.9,-650.8</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>15,-12</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>22,-13.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>15,-15</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>27.5,-13.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>15,-29</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>15,-32</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>10,-11.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>10,-15</position>
<gparam>LABEL_TEXT Input-B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>33.5,-13</position>
<gparam>LABEL_TEXT Output-Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>24,-6.5</position>
<gparam>LABEL_TEXT AND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>22.5,-23</position>
<gparam>LABEL_TEXT OR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>22,-30.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>27.5,-30.5</position>
<input>
<ID>N_in0</ID>7 </input>
<input>
<ID>N_in1</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>10,-28.5</position>
<gparam>LABEL_TEXT Input-A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>10,-31.5</position>
<gparam>LABEL_TEXT Input-B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>33.5,-30</position>
<gparam>LABEL_TEXT Output-Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>22,-37.5</position>
<gparam>LABEL_TEXT NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>BA_NAND2</type>
<position>22,-45</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BE_NOR2</type>
<position>22.5,-58.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>15,-43.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>15,-60</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>15,-57</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>15,-46.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>27.5,-45</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>28,-58.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>22,-52.5</position>
<gparam>LABEL_TEXT NOR gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-14.5,19,-14.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>17 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>17,-15,17,-14.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-12.5,19,-12.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>17 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>17,-12.5,17,-12</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-13.5,26.5,-13.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-29.5,18,-29</points>
<intersection>-29.5 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-29.5,19,-29.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-29,18,-29</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-32,18,-31.5</points>
<intersection>-32 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-31.5,19,-31.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-32,18,-32</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-31.5,27,-31.5</points>
<intersection>26.5 3</intersection>
<intersection>27 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>27,-31.5,27,-31</points>
<intersection>-31.5 1</intersection>
<intersection>-31 7</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-31.5,26.5,-30.5</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>-31.5 1</intersection>
<intersection>-31 7</intersection>
<intersection>-30.5 13</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>26.5,-31,28.5,-31</points>
<intersection>26.5 3</intersection>
<intersection>27 2</intersection>
<intersection>28.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>28.5,-31,28.5,-30.5</points>
<connection>
<GID>26</GID>
<name>N_in1</name></connection>
<intersection>-31 7</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>25,-30.5,26.5,-30.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>26.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-44,18,-43.5</points>
<intersection>-44 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-44,19,-44</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-43.5,18,-43.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-46.5,18,-46</points>
<intersection>-46.5 2</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-46,19,-46</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-46.5,18,-46.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-57.5,19.5,-57.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>18 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-57.5,18,-57</points>
<intersection>-57.5 1</intersection>
<intersection>-57 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,-57,18,-57</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>18 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>19.5,-60,19.5,-59.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-60 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>17,-60,19.5,-60</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>19.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-45,26.5,-45</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-58.5,27,-58.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>50</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>