<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-24.3,12.2667,170.1,-86</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>18,-11.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>11.5,-10.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>11.5,-12.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>22,-11.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>18,-6</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>8.5,-12</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>8.5,-10</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>24.5,-10.5</position>
<gparam>LABEL_TEXT z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>18,-3.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AE_MUX_4x1</type>
<position>17.5,-32</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>11 </output>
<input>
<ID>SEL_0</ID>9 </input>
<input>
<ID>SEL_1</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>12.5,-29</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>12.5,-35</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>12.5,-33</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>12.5,-31</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>19,-25</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>17,-25</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>21.5,-32</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>9.5,-35</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>9.5,-33</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>9.5,-31</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>9.5,-29</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>17,-22.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>19.5,-22.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>24,-31.5</position>
<gparam>LABEL_TEXT z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AI_MUX_8x1</type>
<position>20,-59</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>20 </input>
<input>
<ID>IN_4</ID>19 </input>
<input>
<ID>IN_5</ID>17 </input>
<input>
<ID>IN_6</ID>13 </input>
<input>
<ID>IN_7</ID>12 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>23 </input>
<input>
<ID>SEL_1</ID>22 </input>
<input>
<ID>SEL_2</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>12,-50.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>12,-53</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>12,-65.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>18,-49</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>20,-49</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>22,-49</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>12,-55.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>12,-68</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>12,-60.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>12,-63</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>12,-58</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>24,-59</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>9.5,-67.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>9.5,-65</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>9.5,-62.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>9.5,-60</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>9.5,-57.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>9.5,-55</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>9.5,-52.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>9.5,-50</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>26.5,-58</position>
<gparam>LABEL_TEXT z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>20,-46.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>22.5,-46.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>17.5,-46.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>51.5,-4</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>59,-4</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND3</type>
<position>73,-14.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>38 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND3</type>
<position>73,-22.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>39 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_TOGGLE</type>
<position>67,-4</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND3</type>
<position>73,-30.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<input>
<ID>IN_2</ID>37 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND3</type>
<position>73,-38.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<input>
<ID>IN_2</ID>39 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>77,-14.5</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>77,-22.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>GA_LED</type>
<position>77,-30.5</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>GA_LED</type>
<position>77,-38.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>67,-1.5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>51.5,-1.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>59,-1.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AE_SMALL_INVERTER</type>
<position>54,-9</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_SMALL_INVERTER</type>
<position>62,-9</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>80,-14</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>80,-22</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>80,-30</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>80,-38</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_TOGGLE</type>
<position>105.5,-2</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>113,-2</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>127,-2</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>127,0.5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>105.5,0.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>113,0.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_TOGGLE</type>
<position>120,-2</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>120,0.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AE_SMALL_INVERTER</type>
<position>108,-6</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>AE_SMALL_INVERTER</type>
<position>116,-6</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_SMALL_INVERTER</type>
<position>123,-6</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND4</type>
<position>135,-12</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>53 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND4</type>
<position>135,-22</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>53 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND4</type>
<position>135,-32</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>53 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>139,-12</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>139,-22</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>139,-32</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND4</type>
<position>135,-42</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>53 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>139,-42</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND4</type>
<position>135,-52</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>139,-52</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND4</type>
<position>135,-62</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>52 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>139,-62</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND4</type>
<position>135,-72</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>139,-72</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND4</type>
<position>135,-82</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>58 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>139,-82</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>142.5,-12</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>142,-21.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>142,-32</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>142,-42</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>142,-52</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>142.5,-61.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>142.5,-71.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>142.5,-81.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-10.5,16,-10.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-12.5,16,-12.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-11.5,21,-11.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-9,18,-8</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-29,14.5,-29</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-31,14.5,-31</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-33,14.5,-33</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-35,14.5,-35</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>18.5,-27,19,-27</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>SEL_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-27,17.5,-27</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>SEL_1</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-32,20.5,-32</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<connection>
<GID>19</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-55.5,17,-50.5</points>
<connection>
<GID>42</GID>
<name>IN_7</name></connection>
<intersection>-50.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14,-50.5,17,-50.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-56.5,16.5,-53</points>
<intersection>-56.5 5</intersection>
<intersection>-53 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14,-53,16.5,-53</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>16.5,-56.5,17,-56.5</points>
<connection>
<GID>42</GID>
<name>IN_6</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-65.5,16.5,-65.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>16.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>16.5,-65.5,16.5,-61.5</points>
<intersection>-65.5 1</intersection>
<intersection>-61.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>16.5,-61.5,17,-61.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>16.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-53.5,18,-51</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>18,-53.5,19,-53.5</points>
<connection>
<GID>42</GID>
<name>SEL_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>16,-57.5,16,-55.5</points>
<intersection>-57.5 4</intersection>
<intersection>-55.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-57.5,17,-57.5</points>
<connection>
<GID>42</GID>
<name>IN_5</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>14,-55.5,16,-55.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-68,17,-62.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-68,17,-68</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-58.5,17,-58.5</points>
<connection>
<GID>42</GID>
<name>IN_4</name></connection>
<intersection>13 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>13,-58.5,13,-58</points>
<intersection>-58.5 1</intersection>
<intersection>-58 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>13,-58,14,-58</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>13 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-59.5,17,-59.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>13 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>13,-60.5,13,-59.5</points>
<intersection>-60.5 11</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>13,-60.5,14,-60.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>13 8</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>16,-63,16,-60.5</points>
<intersection>-63 5</intersection>
<intersection>-60.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-60.5,17,-60.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>14,-63,16,-63</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-53.5,20,-51</points>
<connection>
<GID>42</GID>
<name>SEL_1</name></connection>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>22,-53.5,22,-51</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>21,-53.5,22,-53.5</points>
<connection>
<GID>42</GID>
<name>SEL_0</name></connection>
<intersection>22 1</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-59,23,-59</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>42</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-14.5,76,-14.5</points>
<connection>
<GID>101</GID>
<name>N_in0</name></connection>
<connection>
<GID>94</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-22.5,76,-22.5</points>
<connection>
<GID>103</GID>
<name>N_in0</name></connection>
<connection>
<GID>96</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-30.5,76,-30.5</points>
<connection>
<GID>105</GID>
<name>N_in0</name></connection>
<connection>
<GID>98</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-38.5,76,-38.5</points>
<connection>
<GID>107</GID>
<name>N_in0</name></connection>
<connection>
<GID>99</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-32.5,62,-11</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 3</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-14.5,70,-14.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>62,-32.5,70,-32.5</points>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-22.5,54,-11</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 3</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-16.5,70,-16.5</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54,-22.5,70,-22.5</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-40.5,59,-6</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>-40.5 3</intersection>
<intersection>-24.5 1</intersection>
<intersection>-7 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-24.5,70,-24.5</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>59,-40.5,70,-40.5</points>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>59,-7,62,-7</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-38.5,51.5,-6</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 3</intersection>
<intersection>-30.5 1</intersection>
<intersection>-7 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-30.5,70,-30.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>51.5,-38.5,70,-38.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>51.5,-7,54,-7</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-36.5,67,-6</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-36.5 6</intersection>
<intersection>-28.5 7</intersection>
<intersection>-20.5 3</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-12.5,70,-12.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>67,-20.5,70,-20.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>67,-36.5,70,-36.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>67,-28.5,70,-28.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-12,138,-12</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<connection>
<GID>144</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-22,138,-22</points>
<connection>
<GID>150</GID>
<name>N_in0</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-32,138,-32</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<connection>
<GID>146</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-42,138,-42</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<connection>
<GID>153</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-52,138,-52</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<connection>
<GID>155</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-62,138,-62</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<connection>
<GID>157</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-72,138,-72</points>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<connection>
<GID>159</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-82,138,-82</points>
<connection>
<GID>162</GID>
<name>N_in0</name></connection>
<connection>
<GID>161</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-79,127,-4</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>-79 10</intersection>
<intersection>-69 11</intersection>
<intersection>-59 12</intersection>
<intersection>-49 13</intersection>
<intersection>-39 14</intersection>
<intersection>-29 15</intersection>
<intersection>-19 3</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-9,132,-9</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>127,-19,132,-19</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>127,-79,132,-79</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>127,-69,132,-69</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>127,-59,132,-59</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>127,-49,132,-49</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>127,-39,132,-39</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>127,-29,132,-29</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-71,123,-8</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>-71 7</intersection>
<intersection>-51 5</intersection>
<intersection>-31 3</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-11,132,-11</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>123,-31,132,-31</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>123,-51,132,-51</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>123,-71,132,-71</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-63,116,-8</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-63 7</intersection>
<intersection>-53 5</intersection>
<intersection>-23 3</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-13,132,-13</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>116,-23,132,-23</points>
<connection>
<GID>145</GID>
<name>IN_2</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>116,-53,132,-53</points>
<connection>
<GID>155</GID>
<name>IN_2</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>116,-63,132,-63</points>
<connection>
<GID>157</GID>
<name>IN_2</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-45,108,-8</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-45 7</intersection>
<intersection>-35 5</intersection>
<intersection>-25 3</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-15,132,-15</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108,-25,132,-25</points>
<connection>
<GID>145</GID>
<name>IN_3</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>108,-35,132,-35</points>
<connection>
<GID>146</GID>
<name>IN_3</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>108,-45,132,-45</points>
<connection>
<GID>153</GID>
<name>IN_3</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-81,120,-4</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>-81 8</intersection>
<intersection>-61 5</intersection>
<intersection>-41 3</intersection>
<intersection>-21 1</intersection>
<intersection>-4 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-21,132,-21</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>120,-41,132,-41</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>120,-61,132,-61</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>120,-4,123,-4</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>120 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>120,-81,132,-81</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-83,113,-4</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-83 8</intersection>
<intersection>-73 6</intersection>
<intersection>-43 3</intersection>
<intersection>-33 1</intersection>
<intersection>-4 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-33,132,-33</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>113,-43,132,-43</points>
<connection>
<GID>153</GID>
<name>IN_2</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>113,-4,116,-4</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>113,-73,132,-73</points>
<connection>
<GID>159</GID>
<name>IN_2</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>113,-83,132,-83</points>
<connection>
<GID>161</GID>
<name>IN_2</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-85,105.5,-4</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>-85 8</intersection>
<intersection>-75 6</intersection>
<intersection>-65 3</intersection>
<intersection>-55 1</intersection>
<intersection>-4 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-55,132,-55</points>
<connection>
<GID>155</GID>
<name>IN_3</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>105.5,-65,132,-65</points>
<connection>
<GID>157</GID>
<name>IN_3</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>105.5,-4,108,-4</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>105.5,-75,132,-75</points>
<connection>
<GID>159</GID>
<name>IN_3</name></connection>
<intersection>105.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>105.5,-85,132,-85</points>
<connection>
<GID>161</GID>
<name>IN_3</name></connection>
<intersection>105.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>